// Code your testbench here
// or browse Examples

`include "seq_item.sv"
`include "sequence.sv"
`include "sequencer.sv"

`include "driver.sv"
`include "coverage.sv"
`include "monitor.sv"

`include "input_agent.sv"
`include "env.sv"
`include "test.sv"



`include "sap_intf.sv"

`include "top.sv"




